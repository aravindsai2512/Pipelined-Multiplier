// Code your design here
module MULTI_32bit(clk, rst,A, B, F);
   `define BIAS 8'b01111111
   input clk, rst;
   input [31:0]A;
   input [31:0]B;

   output [31:0]F;
   reg [31:0]F;
	

//   reg [1:0]sign;
//   reg [49:0]mantissa;


//////////////// PIPE-LINE REGISTERS /////////////////
reg [62:0] P1;
reg [64:0] P2;
reg [31:0] P3;
//////////////////////////////////////////////////////

initial
begin	
	P1 = 0;
	P2 = 0;
	P3 = 0;
end


wire [1:0]sign;
wire [49:0]mantissa;

assign sign = A[31]+B[31];

//always @ ( F or A or B )
always @ ( posedge clk )
begin
	//solve for the sign bit part
	/////////////////////////////////////////////////////////
	P1[0] <= (sign == 1'b1) ? 1'b1 : 1'b0;
	P1[31:1] <= A[30:0];
	P1[62:32] <= B[30:0];

	///////////////////////////////////////////////////////////
	P2[0] <= P1[0];
	P2[48:1] <={1'b1, P1[23:1]} * {1'b1, P1[54:32]};

	P2[56:49] <= P1[31:24];
	P2[64:57] <= P1[62:55];

///////////////////////////////////////////////////////////
    P3[0] <= P2[0];

    if(P2[48] == 1) begin
	   P3[23:1] = P2[47:25];
       P3[31:24] = P2[56:49] + P2[64:57] - `BIAS + 8'h1;
	end
	else if(P2[47] == 1) begin
	   P3[23:1] = P2[46:24];
       P3[31:24] = P2[56:49] + P2[64:57] - `BIAS ;
	end
	
///////////////////////////////////////////////////////////
	F[31] <= P3[0];
	F[30:0] <= P3[31:1];

////////////////////////////////////////////////////////////
end

endmodule
